library ieee;
use ieee.std_logic_1164.all;

entity tb_gcd  is 
	end tb_gcd;

architecture behavior of tb_gcd is 
signal CLK, RESET: std_logic;
signal A, B, GCD: integer;
component gcd 
	port(CLK, RESET : IN STD_LOGIC;
	    A, B: IN INTEGER;
	    GCD : OUT INTEGER);
END COMPONENT;
BEGIN
gcd1 : gcd port map(CLK=> CLK, RESET=>  RESET, A=>A, B=>B, GCD=>GCD);
clock: process
begin
	CLK<= '1';
	wait for 100 ns;

	CLK <= '0';
	WAIT FOR 100 NS;
	
end process;
process
begin
	RESET <= '1';
	wait for 10 ns;
	RESET  <= '0';

	A <= 10;
	B <= 15;
	wait for 2600 ns;
	
	A <= 3456;
	B <= 234;
	wait for 2600 ns;
	
	A <= 546;
	B <= 24;
	wait for 2600 ns;

	WAIT;
end process;
end behavior;
